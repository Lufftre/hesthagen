library IEEE;
    use IEEE.std_logic_1164.all;
    use IEEE.numeric_std.all;
    use IEEE.std_logic_unsigned.all;
    
entity projectile is
    port (
        CLKPROJECTILE: in std_logic;
        RST: in std_logic;
        pixel_color : out std_logic_vector(2 downto 0)
    );
end entity;

architecture rtl of projectile is 

  signal pixel_counter : integer range 0 to 255 := 0;
  signal rad : std_logic_vector(5 downto 0);
  type projectile_type is array (0 to 255) of std_logic_vector(2 downto 0);
  signal projectile : projectile_type := ("111","111","111","111","111","101","101","101","101","101","101","111","111","111","111","111","111","111","111","101","101","101","101","101","101","101","101","101","101","111","111","111","111","111","101","101","101","101","010","010","010","010","101","101","101","101","111","111","111","101","101","101","010","010","010","010","010","010","010","010","101","101","101","111","111","101","101","010","010","010","010","010","010","010","010","010","010","101","101","111","101","101","101","010","010","010","010","010","010","010","010","010","010","101","101","101","101","101","010","010","010","010","010","010","010","010","010","010","010","010","101","101","101","101","010","010","010","010","010","010","010","010","010","010","010","010","101","101","101","101","010","010","010","010","010","010","010","010","010","010","010","010","101","101","101","101","010","010","010","010","010","010","010","010","010","010","010","010","101","101","101","101","101","010","010","010","010","010","010","010","010","010","010","101","101","101","111","101","101","010","010","010","010","010","010","010","010","010","010","101","101","111","111","101","101","101","010","010","010","010","010","010","010","010","101","101","101","111","111","111","101","101","101","101","010","010","010","010","101","101","101","101","111","111","111","111","111","101","101","101","101","101","101","101","101","101","101","111","111","111","111","111","111","111","111","101","101","101","101","101","101","111","111","111","111","111");

begin 
      -- ----------------------------------------
      --  # Fetching pixelcolor
      -- ----------------------------------------
      process(CLKPROJECTILE) begin
        if rising_edge(CLKPROJECTILE) then
            pixel_color <= projectile(pixel_counter);
            pixel_counter <= pixel_counter + 1;
        end if;
      end process;

end architecture;