library IEEE;
    use IEEE.std_logic_1164.all;
    use IEEE.numeric_std.all;
    use IEEE.std_logic_unsigned.all;
    
entity hest is
    port (
        CLKHORSE: in std_logic;
        RST: in std_logic;
        xctr,yctr : in std_logic_vector(9 downto 0);
        pixel_color : out std_logic_vector(2 downto 0)
    );
end entity;

architecture rtl of hest is 
  signal pixel_counter : std_logic_vector(7 downto 0) := "00000000";
  signal rad : std_logic_vector(5 downto 0);
  type hest_type is array (0 to 255) of std_logic_vector(2 downto 0);
  signal hest : hest_type := (
    "000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000",
    "001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001",
    "000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000",
    "001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001",
    "000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000",
    "001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001",
    "000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000",
    "001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001",
    "000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000",
    "001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001",
    "000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000",
    "001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001",
    "000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000",
    "001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001",
    "000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000",
    "001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"
);

begin 

      -- ----------------------------------------
      --  # Fetching pixelcolor
      -- ----------------------------------------

      process(CLKHORSE) begin
        if rising_edge(CLKHORSE) then
            pixel_color <= hest(conv_integer(pixel_counter));
            pixel_counter <= pixel_counter + 1;
        end if;
      end process;

end architecture;