library IEEE;
    use IEEE.std_logic_1164.all;
    use IEEE.numeric_std.all;
    use IEEE.std_logic_unsigned.all;
    
entity hest is
    port (
        CLKHORSE: in std_logic;
        RST: in std_logic;
        yctr : in integer range 0 to 1023;
        pixel_color : out std_logic_vector(2 downto 0)
    );
end entity;

architecture rtl of hest is 
  signal pixel_counter : integer range 0 to 255 := 0;
  type hest_type is array (0 to 255) of std_logic_vector(2 downto 0);
  signal hest : hest_type := (

"111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","111","111","111","111","111","111","111","111","111","111","111","111","111","000","000","000","000","111","111","111","111","111","111","111","111","111","111","111","000","000","000","000","000","000","000","111","111","111","111","111","111","111","111","111","110","110","110","110","000","000","000","000","111","111","111","111","111","111","111","001","001","110","110","110","110","000","000","000","000","111","111","111","111","111","111","001","110","000","110","110","110","110","000","000","000","000","111","111","111","111","111","001","110","110","110","110","110","110","110","000","000","000","000","111","111","111","001","001","110","110","110","110","110","110","110","110","000","000","000","000","111","111","001","110","110","110","110","110","110","110","110","110","000","000","000","000","111","001","001","110","110","111","111","111","110","110","110","110","000","000","000","000","111","001","110","110","111","111","111","111","110","110","110","110","000","000","000","000","111","001","110","110","111","111","111","111","111","110","110","110","000","000","000","000","111","111","111","111","111","111","111","111","111","110","110","110","000","000","000","000","111","111","111","111","111","111","111","111","111","110","110","110","000","000","000","000","111","111","111","111","111","111","111","111","111","110","110","110","110","110","110","110"

);

begin 

      -- ----------------------------------------
      --  # Fetching pixelcolor
      -- ----------------------------------------

      process(CLKHORSE) begin
        if rising_edge(CLKHORSE) then
            if yctr > 479 - 32 then
              pixel_counter <= 0;
            end if;
            pixel_color <= hest(pixel_counter);
            pixel_counter <= pixel_counter + 1;
        end if;
      end process;

end architecture;