library IEEE;
    use IEEE.std_logic_1164.all;
    use IEEE.numeric_std.all;
    use IEEE.std_logic_unsigned.all;
    
entity hest is
    port (
        CLKHORSE: in std_logic;
        RST: in std_logic;
        xctr,yctr : in std_logic_vector(9 downto 0);
        pixel_color : out std_logic_vector(2 downto 0)
    );
end entity;

architecture rtl of hest is 
  signal pixel_counter : integer range 0 to 255 := 0;
  signal rad : std_logic_vector(5 downto 0);
  type hest_type is array (255 downto to 0) of std_logic_vector(2 downto 0);
  signal hest : hest_type := (

    "000","000","000","000","000","000","000","011","000","000","000","011","000","000","000","000",
    "000","000","000","000","000","000","000","011","000","000","000","011","000","000","000","000",
    "000","000","000","000","100","000","000","011","000","000","000","011","000","000","000","000",
    "000","000","000","000","100","000","000","011","000","000","000","011","000","000","000","000",
    "000","000","000","000","100","000","000","011","000","100","100","011","000","000","000","000",
    "000","000","000","000","000","000","000","011","000","000","000","011","100","000","000","000",
    "000","000","000","000","000","000","000","000","000","000","000","011","000","100","000","000",
    "000","000","000","000","000","000","000","011","000","000","000","011","000","000","000","000",
    "000","000","000","000","000","000","000","011","000","000","000","011","000","000","000","000",
    "000","000","000","000","000","000","000","011","000","000","000","011","000","000","000","000",
    "000","000","000","000","000","000","000","011","000","000","000","011","000","000","000","000",
    "000","000","000","000","000","000","000","011","000","000","000","011","000","000","000","000",
    "000","000","000","000","000","000","000","011","000","000","000","011","000","000","000","000",
    "000","000","000","000","000","000","000","011","000","000","000","011","000","000","000","000",
    "000","000","000","000","000","000","000","011","000","000","000","011","000","000","000","000",
    "000","000","000","000","000","000","000","011","000","000","000","011","000","000","000","000"
);

begin 

      -- ----------------------------------------
      --  # Fetching pixelcolor
      -- ----------------------------------------

      process(CLKHORSE) begin
        if rising_edge(CLKHORSE) then
            pixel_color <= hest(pixel_counter);
            pixel_counter <= pixel_counter + 1;
            if pixel_counter = 255 then
              pixel_counter <= 0;
            end if;
        end if;
      end process;

end architecture;