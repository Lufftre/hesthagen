library IEEE;
    use IEEE.std_logic_1164.all;
    use IEEE.numeric_std.all;
    use IEEE.std_logic_unsigned.all;
    
entity board is
    port (
        CLK: in std_logic;
        RST: in std_logic;
        xctr : in integer range 0 to 1023;
        yctr : in integer range 0 to 1023;
        pixel_color : out std_logic_vector(2 downto 0);
        current_map : in std_logic_vector(2 downto 0)
    );
end entity;

architecture rtl of board is 

  
 signal rad : integer range 0 to 31; 
 signal tile_index : std_logic_vector(11 downto 0);
 signal board_tile : std_logic_vector(1 downto 0);
 signal pixel_color_index : std_logic_vector(2 downto 0);
 signal x : std_logic_vector(9 downto 0);
 signal y : std_logic_vector(9 downto 0);
 

  -- ----------------------------------------
  -- # Colors
  -- ----------------------------------------

  --type colors_type is array (0 to 7) of std_logic_vector(7 downto 0);
  --signal colors : colors_type := (
  --  "000" & "000" & "00", -- BLACK 000
  --  "111" & "111" & "11", -- WHITE 001
  --  "110" & "000" & "00", -- RED   010
  --  "000" & "111" & "00", -- GREEN 011
  --  "000" & "000" & "11", -- BLUE  100
  --  "111" & "000" & "11", -- PINK  101
  --  "000" & "000" & "00", -- MOCHA 110
  --  "100" & "111" & "11" -- ICE    111
  --  );

  --signal colors : colors_type := (
  --  "111" & "111" & "11", -- BLACK 000
  --  "111" & "111" & "11", -- WHITE 001
  --  "000" & "000" & "00", -- RED   010
  --  "111" & "111" & "11", -- GREEN 011
  --  "111" & "111" & "11", -- BLUE  100
  --  "111" & "111" & "11", -- PINK  101
  --  "111" & "111" & "11", -- MOCHA 110
  --  "111" & "111" & "11" -- ICE    111
  --  );
  
  -- ----------------------------------------
  -- # Background tiles
  -- ----------------------------------------

  subtype tmp is std_logic_vector(2 downto 0);
  type tiles_array is array(0 to 3, 0 to 255) of tmp;
  signal pixel_color_array : tiles_array := (

    ("010","010","010","010","010","010","010","101","101","010","010","010","010","010","010","101","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","101","010","010","010","101","010","010","010","010","010","010","010","010","010","010","010","010","010","010","101","101","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","101","101","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","101","010","010","010","101","101","010","010","010","010","010","010","010","010","010","101","010","010","010","010","010","010","010","010","010","101","010","010","101","101","101","010","101","010","010","010","010","010","010","010","010","010","010","010","101","101","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","101","101","101","010","010","010","010","010","010","010","010","010","010","010","010","010","101","010","101","010","010","010","010","010","010","101","010","101","101","010","101","010","010","010","101","010","010","010","010","010","010","010","101","101","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","101","010","010","010","010","010","010","010","010","010","010","010","010","010","010","101","101","010","010","010","010","010","101","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010"),
    ("011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011"),
    ("011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","110","110","110","110","110","110","110","110","110","110","110","110","110","110","011","011","110","110","000","000","000","000","000","000","000","000","000","000","110","110","011","011","110","000","000","110","110","110","110","110","110","110","110","000","000","110","011","011","110","000","110","110","110","110","110","110","110","110","110","110","000","110","011","011","110","000","110","110","110","110","110","110","110","110","110","110","000","110","011","011","110","000","110","110","110","110","110","110","110","110","110","110","000","110","011","011","110","000","110","110","110","110","110","110","110","110","110","110","000","110","011","011","110","000","110","110","110","110","110","110","110","110","110","110","000","110","011","011","110","000","110","110","110","110","110","110","110","110","110","110","000","110","011","011","110","000","110","110","110","110","110","110","110","110","110","110","000","110","011","011","110","000","110","110","110","110","110","110","110","110","110","110","000","110","011","011","110","000","000","110","110","110","110","110","110","110","110","000","000","110","011","011","110","110","000","000","000","000","000","000","000","000","000","000","110","110","011","011","110","110","110","110","110","110","110","110","110","110","110","110","110","110","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011"),
    ("110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","000","000","000","000","000","000","000","000","000","000","110","110","110","110","110","000","000","110","110","110","110","110","110","110","110","000","000","110","110","110","110","000","110","110","110","110","110","110","110","110","110","110","000","110","110","110","110","000","110","110","110","110","110","110","110","110","110","110","000","110","110","110","110","000","110","110","110","110","110","110","110","110","110","110","000","110","110","110","110","000","110","110","110","110","110","110","110","110","110","110","000","110","110","110","110","000","110","110","110","110","110","110","110","110","110","110","000","110","110","110","110","000","110","110","110","110","110","110","110","110","110","110","000","110","110","110","110","000","110","110","110","110","110","110","110","110","110","110","000","110","110","110","110","000","110","110","110","110","110","110","110","110","110","110","000","110","110","110","110","000","000","110","110","110","110","110","110","110","110","000","000","110","110","110","110","110","000","000","000","000","000","000","000","000","000","000","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110")
  );

  
  -- ----------------------------------------
  -- # Board
  -- ----------------------------------------

  type board_type is array (0 to 1023) of std_logic_vector(1 downto 0);

signal board0 : board_type := ("00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","11","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","11","00","00","00","00","00","00","00","00","00","00","00","00","10","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","10","00","00","00","00","00","00","00","00","00","00","00","00","10","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","10","00","00","00","00","00","00","00","00","00","00","00","00","10","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","10","00","00","00","00","00","00","00","00","00","00","00","00","10","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","10","00","00","00","00","00","00","00","00","00","00","00","00","10","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","10","00","00","00","00","00","00","00","00","00","00","00","00","10","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","10","00","00","00","00","00","00","00","00","00","00","00","00","10","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","10","00","00","00","00","00","00","00","00","00","00","00","00","10","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","10","00","00","00","00","00","00","00","00","00","00","00","00","10","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","10","00","00","00","00","00","00","00","00","00","00","00","00","10","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","10","00","00","00","00","00","00","00","00","00","00","00","00","10","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","10","00","00","00","00","00","00","00","00","00","00","00","00","10","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","10","00","00","00","00","00","00","00","00","00","00","00","00","10","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","10","00","00","00","00","00","00","00","00","00","00","00","00","10","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","10","00","00","00","00","00","00","00","00","00","00","00","00","10","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","10","00","00","00","00","00","00","00","00","00","00","00","00","10","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","10","00","00","00","00","00","00","00","00","00","00","00","00","10","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","10","00","00","00","00","00","00","00","00","00","00","00","00","10","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","10","00","00","00","00","00","00","00","00","00","00","00","00","11","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00");
signal board1 : board_type := ("00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","11","10","10","10","10","11","00","00","00","00","00","00","00","00","11","10","10","10","10","11","00","00","00","00","00","00","00","00","00","00","00","00","10","01","01","01","01","10","00","00","00","00","00","00","00","00","10","01","01","01","01","10","00","00","00","00","00","00","00","00","00","00","00","00","10","01","01","01","01","10","00","00","00","00","00","00","00","00","10","01","01","01","01","10","00","00","00","00","00","00","00","00","00","00","00","00","10","01","01","01","01","10","00","00","00","00","00","00","00","00","10","01","01","01","01","10","00","00","00","00","00","00","00","00","00","00","00","00","10","01","01","01","01","10","00","00","00","00","00","00","00","00","10","01","01","01","01","10","00","00","00","00","00","00","00","00","00","00","00","00","11","10","10","10","10","11","00","00","00","00","00","00","00","00","11","10","10","10","10","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","11","10","10","10","10","11","00","00","00","00","00","00","00","00","11","10","10","10","10","11","00","00","00","00","00","00","00","00","00","00","00","00","10","01","01","01","01","10","00","00","00","00","00","00","00","00","10","01","01","01","01","10","00","00","00","00","00","00","00","00","00","00","00","00","10","01","01","01","01","10","00","00","00","00","00","00","00","00","10","01","01","01","01","10","00","00","00","00","00","00","00","00","00","00","00","00","10","01","01","01","01","10","00","00","00","00","00","00","00","00","10","01","01","01","01","10","00","00","00","00","00","00","00","00","00","00","00","00","10","01","01","01","01","10","00","00","00","00","00","00","00","00","10","01","01","01","01","10","00","00","00","00","00","00","00","00","00","00","00","00","11","10","10","10","10","11","00","00","00","00","00","00","00","00","11","10","10","10","10","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00");
signal board2 : board_type := ("00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","11","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","11","00","00","00","00","00","00","00","00","00","00","00","00","10","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","10","00","00","00","00","00","00","00","00","00","00","00","00","10","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","10","00","00","00","00","00","00","00","00","00","00","00","00","10","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","10","00","00","00","00","00","00","00","00","00","00","00","00","10","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","10","00","00","00","00","00","00","00","00","00","00","00","00","10","01","01","01","01","11","10","10","10","10","10","10","10","10","11","01","01","01","01","10","00","00","00","00","00","00","00","00","00","00","00","00","10","01","01","01","01","10","00","00","00","00","00","00","00","00","10","01","01","01","01","10","00","00","00","00","00","00","00","00","00","00","00","00","10","01","01","01","01","10","00","00","00","00","00","00","00","00","10","01","01","01","01","10","00","00","00","00","00","00","00","00","00","00","00","00","10","01","01","01","01","10","00","00","00","00","00","00","00","00","10","01","01","01","01","10","00","00","00","00","00","00","00","00","00","00","00","00","10","01","01","01","01","10","00","00","00","00","00","00","00","00","10","01","01","01","01","10","00","00","00","00","00","00","00","00","00","00","00","00","10","01","01","01","01","10","00","00","00","00","00","00","00","00","10","01","01","01","01","10","00","00","00","00","00","00","00","00","00","00","00","00","10","01","01","01","01","10","00","00","00","00","00","00","00","00","10","01","01","01","01","10","00","00","00","00","00","00","00","00","00","00","00","00","10","01","01","01","01","10","00","00","00","00","00","00","00","00","10","01","01","01","01","10","00","00","00","00","00","00","00","00","00","00","00","00","10","01","01","01","01","10","00","00","00","00","00","00","00","00","10","01","01","01","01","10","00","00","00","00","00","00","00","00","00","00","00","00","10","01","01","01","01","11","10","10","10","10","10","10","10","10","11","01","01","01","01","10","00","00","00","00","00","00","00","00","00","00","00","00","10","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","10","00","00","00","00","00","00","00","00","00","00","00","00","10","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","10","00","00","00","00","00","00","00","00","00","00","00","00","10","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","10","00","00","00","00","00","00","00","00","00","00","00","00","10","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","01","10","00","00","00","00","00","00","00","00","00","00","00","00","11","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","10","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00");
signal board3 : board_type := ("00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","11","10","10","10","10","10","10","10","10","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","10","01","01","01","01","01","01","01","01","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","10","01","01","01","01","01","01","01","01","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","10","01","01","01","01","01","01","01","01","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","10","01","01","01","01","01","01","01","01","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","10","01","01","01","01","01","01","01","01","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","10","01","01","01","01","01","01","01","01","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","10","01","01","01","01","01","01","01","01","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","10","01","01","01","01","01","01","01","01","10","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","11","10","10","10","10","10","10","10","10","11","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00");
signal board4 : board_type := ("00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","01","01","01","01","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","01","00","00","01","00","00","01","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","01","00","00","01","01","00","01","00","00","00","00","00","00","00","01","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","01","01","01","01","00","00","01","00","00","01","01","00","01","00","01","00","00","00","00","00","00","01","01","01","00","00","00","00","00","00","00","00","01","01","00","00","00","00","01","00","01","01","01","01","01","00","01","00","01","01","00","00","01","01","01","01","00","00","00","00","00","00","00","01","01","00","00","00","00","01","01","00","01","01","01","00","01","00","01","01","00","01","00","00","01","01","01","00","01","01","01","00","00","00","00","01","00","00","00","00","00","01","01","00","00","00","00","00","01","00","00","00","01","01","00","00","00","00","00","00","01","01","00","00","00","00","00","01","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","01","01","00","00","00","00","00","00","00","01","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","01","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","01","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","01","00","00","00","01","00","00","00","00","00","00","00","01","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","01","00","00","00","01","01","00","01","00","00","01","00","01","01","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","01","00","00","00","00","01","00","01","00","01","01","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","01","01","00","00","00","00","01","01","01","01","01","00","00","00","00","00","01","00","01","01","01","00","00","01","01","00","00","00","00","00","00","00","01","00","00","00","00","00","01","01","01","01","00","00","00","01","00","00","01","01","01","00","01","01","00","01","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","01","00","00","00","00","01","00","00","01","01","00","00","00","01","00","01","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","01","00","00","00","00","00","00","01","01","00","01","01","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","01","00","00","00","00","00","00","00","00","01","01","01","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00");
signal board5 : board_type := ("00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","01","01","01","00","01","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","01","01","00","01","00","01","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","01","00","01","01","00","01","01","01","01","00","00","01","00","00","00","01","01","01","00","01","00","00","00","00","00","00","00","00","00","00","00","00","01","00","00","00","01","01","01","01","01","01","00","01","00","01","00","01","01","01","00","01","01","01","01","01","01","00","00","00","00","00","00","00","01","00","00","00","01","01","01","01","00","01","00","01","01","01","00","01","00","00","00","01","01","00","00","00","00","00","00","00","00","00","00","00","01","00","00","00","00","00","00","00","00","00","00","00","01","00","00","01","01","01","00","01","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","01","01","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","01","01","01","00","00","00","00","00","00","00","01","01","01","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","01","00","01","01","01","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","01","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","01","01","01","00","00","00","00","01","00","00","00","00","00","00","00","00","00","01","00","00","00","00","00","00","00","00","00","00","00","00","00","01","01","00","00","00","00","00","00","01","00","01","01","00","00","00","01","01","00","01","01","00","00","00","00","00","00","00","00","00","00","00","00","01","00","00","00","00","00","00","00","01","01","01","01","01","01","01","01","00","00","00","01","00","00","00","01","01","00","00","00","00","00","00","00","01","01","01","00","00","00","00","00","01","01","00","00","01","01","00","00","00","00","00","01","00","00","00","01","00","00","00","00","00","00","00","00","00","00","01","01","01","00","00","00","01","01","00","00","01","00","00","00","01","00","00","01","01","01","01","01","01","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","01","00","00","00","00","00","01","00","01","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","01","00","01","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","01","01","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00");

signal current_board : board_type;

begin 
    with current_map select
        current_board <=
            board3 when "000",
            board2 when "001",
            board1 when "010",
            board0 when "011",
            board5 when "101",
            board4 when "110",
        (others => "11") when others;  
      -- ----------------------------------------
      --  # Fetching pixelcolor
      -- ----------------------------------------

      process(CLK) begin
        if rising_edge(CLK) then
            x <= std_logic_vector(to_unsigned(xctr,10));
            y <= std_logic_vector(to_unsigned(yctr,10));
            rad <= yctr/16;
            tile_index <= std_logic_vector(to_unsigned(rad*32 + xctr/16,tile_index'length));

 
            board_tile <= current_board(conv_integer(tile_index));
            pixel_color_index <= pixel_color_array(
                                                  conv_integer(board_tile),
                                                  conv_integer(std_logic_vector((unsigned(y) mod 16)*16) + std_logic_vector((unsigned(x) mod 16)))
                                                  );
            --pixel_color <= colors(conv_integer(pixel_color_index));
            pixel_color <= pixel_color_index;



            --tile_index <= yctr*2 + xctr/16;
            --board_tile <= current_board(tile_index);
            --pixel_color_index <= pixel_color_array(
            --                                      conv_integer(board_tile),
            --                                      (yctr mod 16)*16 + (xctr mod 16)
            --                                      );
            ----pixel_color <= colors(conv_integer(pixel_color_index));
            --pixel_color <= pixel_color_index;

        end if;
      end process;

end architecture;