library IEEE;
    use IEEE.std_logic_1164.all;
    use IEEE.numeric_std.all;
    use IEEE.std_logic_unsigned.all;
    
entity projectile is
    port (
        CLKPROJECTILE: in std_logic;
        RST: in std_logic;
        yctr : in integer range 0 to 1023;
        pixel_color : out std_logic_vector(2 downto 0)
    );
end entity;

architecture rtl of projectile is 

  signal frame_counter : std_logic_vector(5 downto 0) := "000000";
  subtype tmp is std_logic_vector(2 downto 0);
  type frame_array is array(0 to 7, 0 to 255) of tmp;
  signal projectile : frame_array := (


  
  --type projectile_type is array (0 to 255) of std_logic_vector(2 downto 0);
  --signal projectile : projectile_type := 
  ("111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","010","010","010","010","010","010","111","111","111","111","111","111","111","111","010","010","100","100","100","100","100","100","010","010","111","111","111","111","111","111","010","100","101","100","101","100","100","101","100","010","010","111","111","111","111","010","100","101","001","101","101","100","101","101","100","100","010","010","111","111","111","010","100","001","001","101","101","101","101","010","010","010","010","010","010","111","111","010","100","100","001","001","101","100","010","010","111","111","111","010","010","111","111","111","010","100","101","001","101","100","010","111","111","111","111","111","111","111","111","111","010","010","100","100","100","010","010","111","111","111","111","111","111","111","111","111","111","111","010","010","010","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111"),
  ("111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","010","010","111","111","111","111","111","111","111","111","111","111","010","010","010","010","010","010","010","010","111","111","111","111","111","111","111","010","100","010","100","100","010","010","010","111","111","111","111","111","111","111","010","100","100","101","101","100","010","111","111","111","111","111","111","111","111","010","100","100","100","101","101","010","111","111","111","111","111","111","111","111","010","100","100","101","101","101","101","010","111","111","111","111","111","111","111","111","010","100","101","101","101","101","100","100","010","111","111","111","111","111","111","111","010","100","101","101","101","101","101","100","010","111","111","111","111","111","111","111","010","100","101","001","001","001","101","100","010","111","111","111","111","111","111","111","010","100","100","100","100","001","100","010","111","111","111","111","111","111","111","111","010","010","010","010","100","100","010","010","111","111","111","111","111","111","111","111","111","111","111","010","010","010","010","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111"),
  ("111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","010","010","111","111","111","111","111","111","111","111","111","111","111","111","111","010","010","010","111","111","111","111","111","111","111","111","111","111","111","111","010","010","010","111","111","111","111","111","111","111","111","111","111","111","111","010","010","100","010","111","111","111","111","111","111","111","111","111","111","111","111","010","100","100","010","111","111","111","111","111","111","111","111","111","111","111","010","100","101","101","010","010","111","111","111","111","111","111","111","111","111","111","010","100","100","101","101","010","010","010","111","111","111","111","111","111","111","111","010","100","100","100","101","100","100","010","111","111","111","111","111","111","111","111","010","100","101","101","101","101","101","100","010","111","111","111","111","111","111","111","010","100","100","101","101","001","001","100","010","111","111","111","111","111","111","111","010","100","101","001","001","001","101","100","010","111","111","111","111","111","111","111","111","010","100","101","001","100","100","010","111","111","111","111","111","111","111","111","111","010","010","100","100","100","010","010","111","111","111","111","111","111","111","111","111","111","111","010","010","010","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111"),
  ("111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","010","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","010","010","111","111","111","111","111","111","111","111","111","111","111","111","111","010","010","010","111","111","111","111","111","111","111","111","111","111","111","111","111","010","010","010","010","111","111","010","010","010","111","111","111","111","111","111","111","111","010","100","100","010","010","100","100","100","010","010","111","111","111","111","111","111","010","100","101","101","101","100","101","101","100","010","010","111","111","111","111","111","010","010","101","101","101","101","101","001","001","100","010","111","111","111","111","111","010","100","100","100","101","101","101","001","100","100","010","111","111","111","111","111","111","010","100","100","101","101","101","001","100","010","010","111","111","111","111","111","111","111","010","100","100","101","101","101","100","010","111","111","111","111","111","111","111","111","111","010","100","100","100","100","100","010","111","111","111","111","111","111","111","111","111","111","010","010","010","010","010","010","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111"),
  ("111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","010","010","010","111","111","111","111","111","111","111","111","111","111","111","010","010","100","100","100","010","010","111","111","111","111","111","111","111","111","111","010","100","101","001","101","100","010","111","111","111","010","010","111","111","111","010","010","100","101","001","001","100","100","010","111","111","010","010","010","010","010","010","101","101","101","101","001","001","100","010","111","111","111","010","010","100","100","101","101","100","101","101","001","101","100","010","111","111","111","111","010","010","100","101","100","100","101","100","101","100","010","111","111","111","111","111","111","010","010","100","100","100","100","100","100","010","010","111","111","111","111","111","111","111","111","010","010","010","010","010","010","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111"),
  ("111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","010","010","010","010","111","111","111","111","111","111","111","111","111","111","111","010","010","100","100","010","010","010","010","111","111","111","111","111","111","111","111","010","100","001","100","100","100","100","010","111","111","111","111","111","111","111","010","100","101","001","001","001","101","100","010","111","111","111","111","111","111","111","010","100","101","101","101","101","101","100","010","111","111","111","111","111","111","111","010","100","100","101","101","101","101","100","010","111","111","111","111","111","111","111","111","010","101","101","101","101","100","100","010","111","111","111","111","111","111","111","111","010","101","101","100","100","100","010","111","111","111","111","111","111","111","111","010","100","101","101","100","100","010","111","111","111","111","111","111","111","010","010","010","100","100","010","100","010","111","111","111","111","111","111","111","010","010","010","010","010","010","010","010","111","111","111","111","111","111","111","111","111","111","010","010","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111"),
  ("111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","010","010","010","111","111","111","111","111","111","111","111","111","111","111","010","010","100","100","100","010","010","111","111","111","111","111","111","111","111","111","010","100","100","001","101","100","010","111","111","111","111","111","111","111","111","010","100","101","001","001","001","101","100","010","111","111","111","111","111","111","111","010","100","001","001","101","101","100","100","010","111","111","111","111","111","111","111","010","100","101","101","101","101","101","100","010","111","111","111","111","111","111","111","111","010","100","100","101","100","100","100","010","111","111","111","111","111","111","111","111","010","010","010","101","101","100","100","010","111","111","111","111","111","111","111","111","111","111","010","010","101","101","100","010","111","111","111","111","111","111","111","111","111","111","111","010","100","100","010","111","111","111","111","111","111","111","111","111","111","111","111","010","100","010","010","111","111","111","111","111","111","111","111","111","111","111","111","010","010","010","111","111","111","111","111","111","111","111","111","111","111","111","010","010","010","111","111","111","111","111","111","111","111","111","111","111","111","111","010","010","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111"),
  ("111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","010","010","010","010","111","111","111","111","111","111","111","111","111","111","111","010","100","100","100","100","010","111","111","111","111","111","111","111","111","111","010","010","100","101","101","100","100","010","111","111","111","111","111","111","111","111","010","100","001","101","101","100","100","100","010","111","111","111","111","111","111","010","010","100","001","001","101","101","101","100","100","010","111","111","111","111","111","111","010","100","001","001","101","101","100","100","100","010","111","111","111","111","111","111","010","100","001","101","100","101","100","101","101","010","010","111","111","111","111","111","010","010","100","101","010","010","101","101","100","010","010","111","111","111","111","111","111","010","010","010","010","111","010","010","100","010","010","111","111","111","111","111","111","111","111","111","111","111","111","111","010","010","010","111","111","111","111","111","111","111","111","111","111","111","111","111","111","010","010","111","111","111","111","111","111","111","111","111","111","111","111","111","111","010","010","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111")
  
  );
  signal pixel_counter : integer range 0 to 255 := 1;
begin 
      -- ----------------------------------------
      --  # Fetching pixelcolor
      -- ----------------------------------------
      process(CLKPROJECTILE) begin
        if rising_edge(CLKPROJECTILE) then
            if yctr > 479 - 32 then
              pixel_counter <= 0;
            end if;
            if pixel_counter = 255 then
              frame_counter <= frame_counter + 1;
            end if;
            pixel_color <= projectile(conv_integer(frame_counter(5 downto 3)),pixel_counter);
            pixel_counter <= pixel_counter + 1;
        end if;
      end process;

end architecture;